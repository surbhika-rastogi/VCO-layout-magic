magic
tech min2
timestamp 1465277592
<< nwell >>
rect -1 0 25 27
<< ntransistor >>
rect 11 -16 13 -6
<< ptransistor >>
rect 11 6 13 16
<< ndiffusion >>
rect 10 -16 11 -6
rect 13 -16 14 -6
<< pdiffusion >>
rect 10 6 11 16
rect 13 6 14 16
<< ndcontact >>
rect 6 -16 10 -6
rect 14 -16 18 -6
<< pdcontact >>
rect 6 6 10 16
rect 14 6 18 16
<< psubstratepcontact >>
rect 2 -28 6 -24
rect 10 -28 14 -24
rect 18 -28 22 -24
<< nsubstratencontact >>
rect 2 20 6 24
rect 10 20 14 24
rect 18 20 22 24
<< polysilicon >>
rect 11 16 13 19
rect 11 -2 13 6
rect 3 -4 13 -2
rect 11 -6 13 -4
rect 11 -19 13 -16
<< polycontact >>
rect -1 -5 3 -1
<< metal1 >>
rect 0 20 2 24
rect 6 16 10 24
rect 14 20 18 24
rect 22 20 24 24
rect 14 -1 18 6
rect -3 -5 -1 -1
rect 14 -5 22 -1
rect 14 -6 18 -5
rect 6 -28 10 -16
rect 14 -28 18 -24
<< labels >>
rlabel metal1 23 21 23 21 7 vdd!
rlabel metal1 -3 -5 -3 -1 3 in
rlabel metal1 22 -5 22 -1 7 out
rlabel metal1 15 -27 15 -27 1 gnd!
<< end >>
